module mux4( select, d, q );

input[1:0] select;
input[9:0] d[3:0];
output [9:0] q;

reg       q;
wire[1:0] select;
wire[3:0] d;

always @( select or d )
begin
   case( select )
       0 : q = d[0];
       1 : q = d[1];
       2 : q = d[2];
       3 : q = d[3];
   endcase
end

endmodule
